module adder_para
    # (parameter N=4)
    (
        input wire [N-1:0] a,b,
        output reg [N-1:0] sum,
        output reg cout
    );
    localparam N1 = N-1;
    assign var = value;
endmodule
